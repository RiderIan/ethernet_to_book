`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Ian Rider
// 
//////////////////////////////////////////////////////////////////////////////////

module RGMII_TX (
    input  logic rstIn,
    input  logic clk125In,
    input  logic intBIn,

    output logic txDataOut,
    output logic txCtrlOut);

endmodule